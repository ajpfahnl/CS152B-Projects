module alu16

endmodule