module alu16(A, B, ALUCtrl, S, Zero, Overflow);
    input wire [15:0] A, B,
    wire [3:0] ALUCtrl,
    output wire [15:0] S,
    Zero, Overflow;

    // run all ALU operations
    mux161()
endmodule